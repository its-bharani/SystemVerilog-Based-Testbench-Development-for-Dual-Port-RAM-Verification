interface ram_if(input bit clk);
  logic [
